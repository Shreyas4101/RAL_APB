// FRONTDOOR

`include "sequences/fctrl_seq.sv"
`include "sequences/fr1_seq.sv"
`include "sequences/fr2_seq.sv"
`include "sequences/fr3_seq.sv"
`include "sequences/fr4_seq.sv"
//`include "sequences/freg_seq.sv"
`include "sequences/rst1_seq.sv"
`include "sequences/rst2_seq.sv"
`include "sequences/rst3_seq.sv"
`include "sequences/rst4_seq.sv"
