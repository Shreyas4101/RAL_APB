`include "sequences/br1_seq.sv"
`include "sequences/br2_seq.sv"
`include "sequences/br3_seq.sv"
`include "sequences/br4_seq.sv"
`include "sequences/bctrl_seq.sv"
