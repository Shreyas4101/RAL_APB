// FRONTDOOR

`include "sequences/frontdoor/fr1_seq.sv"
`include "sequences/frontdoor/fr2_seq.sv"
`include "sequences/frontdoor/fr3_seq.sv"
`include "sequences/frontdoor/fr4_seq.sv"
//`include "sequences/frontdoor/freg_seq.sv"
`include "sequences/frontdoor/rst1_seq.sv"
`include "sequences/frontdoor/rst2_seq.sv"
`include "sequences/frontdoor/rst3_seq.sv"
`include "sequences/frontdoor/rst4_seq.sv"


// BACKDOOR

`include "sequences/backdoor/br1_seq.sv"
`include "sequences/backdoor/br2_seq.sv"
`include "sequences/backdoor/br3_seq.sv"
`include "sequences/backdoor/br4_seq.sv"
//`include "sequences/backdoor/breg_seq.sv"
