`include "ral_interface.sv"
`include "ral_reg.sv"
`include "ral_regblock.sv"
`include "ral_seq_item.sv"
`include "ral_adapter.sv"
`include "ral_reg_seq.sv"
//`include "sequence.sv"
`include "ral_sequencer.sv"
`include "ral_driver.sv"
`include "ral_monitor.sv"
`include "ral_agent.sv"
`include "ral_scb.sv"
`include "ral_env.sv"
`include "ral_test.sv"
